TCM_AHBL_Adapter.FSM.bsv